`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/08/2021 05:21:11 AM
// Design Name: 
// Module Name: pipeline_sort
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`default_nettype none
module pipeline_sort(
        input wire clk, 
        input wire rst, 
        input wire start, 
        output logic done_out
        
         
    );
endmodule
`default_nettype wire
